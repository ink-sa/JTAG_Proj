`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:39:36 12/23/2016 
// Design Name: 
// Module Name:    BIST_mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BIST_mem #(parameter N = 8, M = 16) //2^8 ����� ������ �� 16 ��� ������
   (input clk,
    input we,
    input res,
    input [N-1:0] adr,
    input [M-1:0] in,
    output [M-1:0] out
    );
	
	reg [M-1:0] mem [2**N-1:0];
	
	integer i;
	
	always @(posedge clk) begin
		if (res) begin						
		//������������� ������
				mem [0] <= 16'h20_00;
				mem [1] <= 16'h12_01;
				mem [2] <= 16'h1A_13;
				mem [3] <= 16'h1A_34;
				mem [4] <= 16'h1F_41;
				mem [5] <= 16'h20_00;
				mem [6] <= 16'h12_01;
				mem [7] <= 16'h1A_13;
				mem [8] <= 16'h1A_34;
				mem [9] <= 16'h11_47;
				mem [10] <= 16'h20_00;
				mem [11] <= 16'h12_01;
				mem [12] <= 16'h1A_13;
				mem [13] <= 16'h1A_34;
				mem [14] <= 16'h1E_49;
				mem [15] <= 16'h20_00;
				mem [16] <= 16'h12_01;
				mem [17] <= 16'h1A_13;
				mem [18] <= 16'h1A_34;
				mem [19] <= 16'h15_4C;
				mem [20] <= 16'h20_00;
				mem [21] <= 16'h12_01;
				mem [22] <= 16'h12_1B;
				mem [23] <= 16'h1D_B8;
				mem [24] <= 16'h1D_83;
				mem [25] <= 16'h20_00;
				mem [26] <= 16'h12_01;
				mem [27] <= 16'h12_1B;
				mem [28] <= 16'h1D_B8;
				mem [29] <= 16'h13_87;
				mem [30] <= 16'h20_00;
				mem [31] <= 16'h12_01;
				mem [32] <= 16'h12_1B;
				mem [33] <= 16'h1D_B8;
				mem [34] <= 16'h1F_8B;
				mem [35] <= 16'h20_00;
				mem [36] <= 16'h12_01;
				mem [37] <= 16'h12_1B;
				mem [38] <= 16'h19_BE;
				mem [39] <= 16'h1F_E1;
				mem [40] <= 16'h20_00;
				mem [41] <= 16'h12_01;
				mem [42] <= 16'h12_1B;
				mem [43] <= 16'h19_BE;
				mem [44] <= 16'h1D_E4;
				mem [45] <= 16'h20_00;
				mem [46] <= 16'h12_01;
				mem [47] <= 16'h12_1B;
				mem [48] <= 16'h19_BE;
				mem [49] <= 16'h1C_E7;
				mem [50] <= 16'h20_00;
				mem [51] <= 16'h18_06;
				mem [52] <= 16'h13_69;
				mem [53] <= 16'h11_97;
				mem [54] <= 16'h10_70;
				mem [55] <= 16'h20_00;
				mem [56] <= 16'h18_06;
				mem [57] <= 16'h13_69;
				mem [58] <= 16'h11_97;
				mem [59] <= 16'h1E_72;
				mem [60] <= 16'h20_00;
				mem [61] <= 16'h18_06;
				mem [62] <= 16'h13_69;
				mem [63] <= 16'h11_97;
				mem [64] <= 16'h15_75;
				mem [65] <= 16'h20_00;
				mem [66] <= 16'h18_06;
				mem [67] <= 16'h13_69;
				mem [68] <= 16'h11_97;
				mem [69] <= 16'h13_7A;
				mem [70] <= 16'h20_00;
				mem [71] <= 16'h18_06;
				mem [72] <= 16'h13_69;
				mem [73] <= 16'h11_97;
				mem [74] <= 16'h1F_7E;
				mem [75] <= 16'h20_00;
				mem [76] <= 16'h1F_0D;
				mem [77] <= 16'h17_DF;
				mem [78] <= 16'h10_FA;
				mem [79] <= 16'h13_A2;
				mem [80] <= 16'h20_00;
				mem [81] <= 16'h1F_0D;
				mem [82] <= 16'h17_DF;
				mem [83] <= 16'h10_FA;
				mem [84] <= 16'h1F_A5;
				mem [85] <= 16'h20_00;
				mem [86] <= 16'h1F_0D;
				mem [87] <= 16'h17_DF;
				mem [88] <= 16'h10_FA;
				mem [89] <= 16'h1A_A8;
				mem [90] <= 16'h20_00;
				mem [91] <= 16'h1F_0D;
				mem [92] <= 16'h17_DF;
				mem [93] <= 16'h10_FA;
				mem [94] <= 16'h11_AD;
				mem [95] <= 16'h20_00;
				mem [96] <= 16'h12_01;
				mem [97] <= 16'h1A_13;
				mem [98] <= 16'h1E_32;
				mem [99] <= 16'h20_00;
				mem [100] <= 16'h12_01;
				mem [101] <= 16'h1A_13;
				mem [102] <= 16'h1A_34;
				mem [103] <= 16'h20_00;
				mem [104] <= 16'h12_01;
				mem [105] <= 16'h1A_13;
				mem [106] <= 16'h16_3D;
				mem [107] <= 16'h20_00;
				mem [108] <= 16'h12_01;
				mem [109] <= 16'h12_1B;
				mem [110] <= 16'h1A_B1;
				mem [111] <= 16'h20_00;
				mem [112] <= 16'h12_01;
				mem [113] <= 16'h12_1B;
				mem [114] <= 16'h1D_B8;
				mem [115] <= 16'h20_00;
				mem [116] <= 16'h12_01;
				mem [117] <= 16'h12_1B;
				mem [118] <= 16'h1E_BC;
				mem [119] <= 16'h20_00;
				mem [120] <= 16'h12_01;
				mem [121] <= 16'h12_1B;
				mem [122] <= 16'h19_BE;
				mem [123] <= 16'h20_00;
				mem [124] <= 16'h18_06;
				mem [125] <= 16'h10_62;
				mem [126] <= 16'h1B_21;
				mem [127] <= 16'h20_00;
				mem [128] <= 16'h18_06;
				mem [129] <= 16'h10_62;
				mem [130] <= 16'h1F_26;
				mem [131] <= 16'h20_00;
				mem [132] <= 16'h18_06;
				mem [133] <= 16'h10_62;
				mem [134] <= 16'h10_29;
				mem [135] <= 16'h20_00;
				mem [136] <= 16'h18_06;
				mem [137] <= 16'h10_62;
				mem [138] <= 16'h1C_2E;
				mem [139] <= 16'h20_00;
				mem [140] <= 16'h18_06;
				mem [141] <= 16'h11_65;
				mem [142] <= 16'h1C_50;
				mem [143] <= 16'h20_00;
				mem [144] <= 16'h18_06;
				mem [145] <= 16'h11_65;
				mem [146] <= 16'h13_52;
				mem [147] <= 16'h20_00;
				mem [148] <= 16'h18_06;
				mem [149] <= 16'h11_65;
				mem [150] <= 16'h1F_54;
				mem [151] <= 16'h20_00;
				mem [152] <= 16'h18_06;
				mem [153] <= 16'h11_65;
				mem [154] <= 16'h12_58;
				mem [155] <= 16'h20_00;
				mem [156] <= 16'h18_06;
				mem [157] <= 16'h11_65;
				mem [158] <= 16'h1D_5D;
				mem [159] <= 16'h20_00;
				mem [160] <= 16'h18_06;
				mem [161] <= 16'h13_69;
				mem [162] <= 16'h10_94;
				mem [163] <= 16'h20_00;
				mem [164] <= 16'h18_06;
				mem [165] <= 16'h13_69;
				mem [166] <= 16'h11_97;
				mem [167] <= 16'h20_00;
				mem [168] <= 16'h18_06;
				mem [169] <= 16'h13_69;
				mem [170] <= 16'h1E_9C;
				mem [171] <= 16'h20_00;
				mem [172] <= 16'h18_06;
				mem [173] <= 16'h13_69;
				mem [174] <= 16'h1B_9E;
				mem [175] <= 16'h20_00;
				mem [176] <= 16'h18_06;
				mem [177] <= 16'h1F_6C;
				mem [178] <= 16'h1E_C3;
				mem [179] <= 16'h20_00;
				mem [180] <= 16'h18_06;
				mem [181] <= 16'h1F_6C;
				mem [182] <= 16'h19_C6;
				mem [183] <= 16'h20_00;
				mem [184] <= 16'h18_06;
				mem [185] <= 16'h1F_6C;
				mem [186] <= 16'h1B_C9;
				mem [187] <= 16'h20_00;
				mem [188] <= 16'h18_06;
				mem [189] <= 16'h1F_6C;
				mem [190] <= 16'h12_CE;
				mem [191] <= 16'h20_00;
				mem [192] <= 16'h1F_0D;
				mem [193] <= 16'h17_DF;
				mem [194] <= 16'h1C_F3;
				mem [195] <= 16'h20_00;
				mem [196] <= 16'h1F_0D;
				mem [197] <= 16'h17_DF;
				mem [198] <= 16'h1A_F7;
				mem [199] <= 16'h20_00;
				mem [200] <= 16'h1F_0D;
				mem [201] <= 16'h17_DF;
				mem [202] <= 16'h10_FA;
				mem [203] <= 16'h20_00;
				mem [204] <= 16'h1F_0D;
				mem [205] <= 16'h17_DF;
				mem [206] <= 16'h14_FC;
				mem [207] <= 16'h20_00;
				mem [208] <= 16'h12_01;
				mem [209] <= 16'h17_10;
				mem [210] <= 16'h20_00;
				mem [211] <= 16'h12_01;
				mem [212] <= 16'h1A_13;
				mem [213] <= 16'h20_00;
				mem [214] <= 16'h12_01;
				mem [215] <= 16'h12_1B;
				mem [216] <= 16'h20_00;
				mem [217] <= 16'h18_06;
				mem [218] <= 16'h10_62;
				mem [219] <= 16'h20_00;
				mem [220] <= 16'h18_06;
				mem [221] <= 16'h11_65;
				mem [222] <= 16'h20_00;
				mem [223] <= 16'h18_06;
				mem [224] <= 16'h13_69;
				mem [225] <= 16'h20_00;
				mem [226] <= 16'h18_06;
				mem [227] <= 16'h1F_6C;
				mem [228] <= 16'h20_00;
				mem [229] <= 16'h1F_0D;
				mem [230] <= 16'h15_D2;
				mem [231] <= 16'h20_00;
				mem [232] <= 16'h1F_0D;
				mem [233] <= 16'h19_D3;
				mem [234] <= 16'h20_00;
				mem [235] <= 16'h1F_0D;
				mem [236] <= 16'h1E_D5;
				mem [237] <= 16'h20_00;
				mem [238] <= 16'h1F_0D;
				mem [239] <= 16'h1F_D9;
				mem [240] <= 16'h20_00;
				mem [241] <= 16'h1F_0D;
				mem [242] <= 16'h17_DF; 
				mem [243] <= 16'h20_00;

				for(i=244; i < 2**N; i = i + 1) begin
					mem[i] <= 16'h0000;						//����������� ����������� ������ BIST �� ������/���������
				end				
		end
		else if (we) mem[adr] <= in;
	end
	assign out = mem[adr];

endmodule
